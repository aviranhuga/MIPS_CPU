
LIBRARY IEEE; 		
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY WRITEBACK IS
	  PORT(	
			read_data 	: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			ALU_result	: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			MemtoReg    : IN    STD_LOGIC;
			write_data 	: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 ));
END WRITEBACK;

ARCHITECTURE behavior OF WRITEBACK IS

BEGIN
	write_data <= ALU_result( 31 DOWNTO 0 ) 
			WHEN ( MemtoReg = '0' ) 	ELSE read_data;
		
END behavior;


